magic
tech sky130A
magscale 1 2
timestamp 1702659099
<< nwell >>
rect 760 2352 1212 3590
rect 1600 2339 2052 3577
rect 2479 2414 2931 3652
rect 3319 2401 3771 3639
rect 750 800 1232 2038
rect 1610 790 2092 2028
rect 2450 810 2932 2048
rect 3270 800 3752 2038
<< pwell >>
rect -4115 57 -4049 109
rect 757 -43 1239 777
rect 1617 -53 2099 767
rect 2457 -33 2939 787
rect 3277 -43 3759 777
rect 780 -1390 1232 -170
rect 1650 -1370 2102 -150
rect 2480 -1380 2932 -160
rect 3290 -1360 3742 -140
<< nmos >>
rect 953 167 1043 567
rect 1813 157 1903 557
rect 2653 177 2743 577
rect 3473 167 3563 567
rect 976 -1180 1036 -380
rect 1846 -1160 1906 -360
rect 2676 -1170 2736 -370
rect 3486 -1150 3546 -350
<< pmos >>
rect 956 2571 1016 3371
rect 1796 2558 1856 3358
rect 2675 2633 2735 3433
rect 3515 2620 3575 3420
rect 946 1019 1036 1819
rect 1806 1009 1896 1809
rect 2646 1029 2736 1829
rect 3466 1019 3556 1819
<< ndiff >>
rect 895 555 953 567
rect 895 179 907 555
rect 941 179 953 555
rect 895 167 953 179
rect 1043 555 1101 567
rect 1043 179 1055 555
rect 1089 179 1101 555
rect 1043 167 1101 179
rect 1755 545 1813 557
rect 1755 169 1767 545
rect 1801 169 1813 545
rect 1755 157 1813 169
rect 1903 545 1961 557
rect 1903 169 1915 545
rect 1949 169 1961 545
rect 1903 157 1961 169
rect 2595 565 2653 577
rect 2595 189 2607 565
rect 2641 189 2653 565
rect 2595 177 2653 189
rect 2743 565 2801 577
rect 2743 189 2755 565
rect 2789 189 2801 565
rect 2743 177 2801 189
rect 3415 555 3473 567
rect 3415 179 3427 555
rect 3461 179 3473 555
rect 3415 167 3473 179
rect 3563 555 3621 567
rect 3563 179 3575 555
rect 3609 179 3621 555
rect 3563 167 3621 179
rect 918 -392 976 -380
rect 918 -1168 930 -392
rect 964 -1168 976 -392
rect 918 -1180 976 -1168
rect 1036 -392 1094 -380
rect 1036 -1168 1048 -392
rect 1082 -1168 1094 -392
rect 1036 -1180 1094 -1168
rect 1788 -372 1846 -360
rect 1788 -1148 1800 -372
rect 1834 -1148 1846 -372
rect 1788 -1160 1846 -1148
rect 1906 -372 1964 -360
rect 1906 -1148 1918 -372
rect 1952 -1148 1964 -372
rect 1906 -1160 1964 -1148
rect 2618 -382 2676 -370
rect 2618 -1158 2630 -382
rect 2664 -1158 2676 -382
rect 2618 -1170 2676 -1158
rect 2736 -382 2794 -370
rect 2736 -1158 2748 -382
rect 2782 -1158 2794 -382
rect 2736 -1170 2794 -1158
rect 3428 -362 3486 -350
rect 3428 -1138 3440 -362
rect 3474 -1138 3486 -362
rect 3428 -1150 3486 -1138
rect 3546 -362 3604 -350
rect 3546 -1138 3558 -362
rect 3592 -1138 3604 -362
rect 3546 -1150 3604 -1138
<< pdiff >>
rect 898 3359 956 3371
rect 898 2583 910 3359
rect 944 2583 956 3359
rect 898 2571 956 2583
rect 1016 3359 1074 3371
rect 1016 2583 1028 3359
rect 1062 2583 1074 3359
rect 1016 2571 1074 2583
rect 1738 3346 1796 3358
rect 1738 2570 1750 3346
rect 1784 2570 1796 3346
rect 1738 2558 1796 2570
rect 1856 3346 1914 3358
rect 1856 2570 1868 3346
rect 1902 2570 1914 3346
rect 1856 2558 1914 2570
rect 2617 3421 2675 3433
rect 2617 2645 2629 3421
rect 2663 2645 2675 3421
rect 2617 2633 2675 2645
rect 2735 3421 2793 3433
rect 2735 2645 2747 3421
rect 2781 2645 2793 3421
rect 2735 2633 2793 2645
rect 3457 3408 3515 3420
rect 3457 2632 3469 3408
rect 3503 2632 3515 3408
rect 3457 2620 3515 2632
rect 3575 3408 3633 3420
rect 3575 2632 3587 3408
rect 3621 2632 3633 3408
rect 3575 2620 3633 2632
rect 888 1807 946 1819
rect 888 1031 900 1807
rect 934 1031 946 1807
rect 888 1019 946 1031
rect 1036 1807 1094 1819
rect 1036 1031 1048 1807
rect 1082 1031 1094 1807
rect 1036 1019 1094 1031
rect 1748 1797 1806 1809
rect 1748 1021 1760 1797
rect 1794 1021 1806 1797
rect 1748 1009 1806 1021
rect 1896 1797 1954 1809
rect 1896 1021 1908 1797
rect 1942 1021 1954 1797
rect 1896 1009 1954 1021
rect 2588 1817 2646 1829
rect 2588 1041 2600 1817
rect 2634 1041 2646 1817
rect 2588 1029 2646 1041
rect 2736 1817 2794 1829
rect 2736 1041 2748 1817
rect 2782 1041 2794 1817
rect 2736 1029 2794 1041
rect 3408 1807 3466 1819
rect 3408 1031 3420 1807
rect 3454 1031 3466 1807
rect 3408 1019 3466 1031
rect 3556 1807 3614 1819
rect 3556 1031 3568 1807
rect 3602 1031 3614 1807
rect 3556 1019 3614 1031
<< ndiffc >>
rect 907 179 941 555
rect 1055 179 1089 555
rect 1767 169 1801 545
rect 1915 169 1949 545
rect 2607 189 2641 565
rect 2755 189 2789 565
rect 3427 179 3461 555
rect 3575 179 3609 555
rect 930 -1168 964 -392
rect 1048 -1168 1082 -392
rect 1800 -1148 1834 -372
rect 1918 -1148 1952 -372
rect 2630 -1158 2664 -382
rect 2748 -1158 2782 -382
rect 3440 -1138 3474 -362
rect 3558 -1138 3592 -362
<< pdiffc >>
rect 910 2583 944 3359
rect 1028 2583 1062 3359
rect 1750 2570 1784 3346
rect 1868 2570 1902 3346
rect 2629 2645 2663 3421
rect 2747 2645 2781 3421
rect 3469 2632 3503 3408
rect 3587 2632 3621 3408
rect 900 1031 934 1807
rect 1048 1031 1082 1807
rect 1760 1021 1794 1797
rect 1908 1021 1942 1797
rect 2600 1041 2634 1817
rect 2748 1041 2782 1817
rect 3420 1031 3454 1807
rect 3568 1031 3602 1807
<< psubdiff >>
rect 793 707 1203 741
rect 793 645 827 707
rect 793 27 827 89
rect 1169 27 1203 707
rect 793 -7 1203 27
rect 1653 697 2063 731
rect 1653 635 1687 697
rect 1653 17 1687 79
rect 2029 17 2063 697
rect 1653 -17 2063 17
rect 2493 717 2903 751
rect 2493 655 2527 717
rect 2493 37 2527 99
rect 2869 37 2903 717
rect 2493 3 2903 37
rect 3313 707 3723 741
rect 3313 645 3347 707
rect 3313 27 3347 89
rect 3689 27 3723 707
rect 3313 -7 3723 27
rect 816 -240 1196 -206
rect 816 -1320 850 -240
rect 1162 -1320 1196 -240
rect 816 -1354 912 -1320
rect 1100 -1354 1196 -1320
rect 1686 -220 2066 -186
rect 1686 -1300 1720 -220
rect 2032 -1300 2066 -220
rect 1686 -1334 1782 -1300
rect 1970 -1334 2066 -1300
rect 2516 -230 2896 -196
rect 2516 -1310 2550 -230
rect 2862 -1310 2896 -230
rect 2516 -1344 2612 -1310
rect 2800 -1344 2896 -1310
rect 3326 -210 3706 -176
rect 3326 -1290 3360 -210
rect 3672 -1290 3706 -210
rect 3326 -1324 3422 -1290
rect 3610 -1324 3706 -1290
<< nsubdiff >>
rect 2515 3582 2611 3616
rect 2799 3582 2895 3616
rect 796 3520 892 3554
rect 1080 3520 1176 3554
rect 796 2422 830 3520
rect 1142 2422 1176 3520
rect 796 2388 1176 2422
rect 1636 3507 1732 3541
rect 1920 3507 2016 3541
rect 1636 2409 1670 3507
rect 1982 2409 2016 3507
rect 2515 2484 2549 3582
rect 2861 2484 2895 3582
rect 2515 2450 2895 2484
rect 3355 3569 3451 3603
rect 3639 3569 3735 3603
rect 3355 2471 3389 3569
rect 3701 2471 3735 3569
rect 3355 2437 3735 2471
rect 1636 2375 2016 2409
rect 786 1968 1196 2002
rect 786 1906 820 1968
rect 786 870 820 932
rect 1162 870 1196 1968
rect 786 836 1196 870
rect 1646 1958 2056 1992
rect 1646 1896 1680 1958
rect 1646 860 1680 922
rect 2022 860 2056 1958
rect 1646 826 2056 860
rect 2486 1978 2896 2012
rect 2486 1916 2520 1978
rect 2486 880 2520 942
rect 2862 880 2896 1978
rect 2486 846 2896 880
rect 3306 1968 3716 2002
rect 3306 1906 3340 1968
rect 3306 870 3340 932
rect 3682 870 3716 1968
rect 3306 836 3716 870
<< psubdiffcont >>
rect 793 89 827 645
rect 1653 79 1687 635
rect 2493 99 2527 655
rect 3313 89 3347 645
rect 912 -1354 1100 -1320
rect 1782 -1334 1970 -1300
rect 2612 -1344 2800 -1310
rect 3422 -1324 3610 -1290
<< nsubdiffcont >>
rect 2611 3582 2799 3616
rect 892 3520 1080 3554
rect 1732 3507 1920 3541
rect 3451 3569 3639 3603
rect 786 932 820 1906
rect 1646 922 1680 1896
rect 2486 942 2520 1916
rect 3306 932 3340 1906
<< poly >>
rect 953 3452 1019 3468
rect 953 3418 969 3452
rect 1003 3418 1019 3452
rect 953 3402 1019 3418
rect 956 3371 1016 3402
rect 956 2540 1016 2571
rect 953 2524 1019 2540
rect 953 2490 969 2524
rect 1003 2490 1019 2524
rect 953 2474 1019 2490
rect 1793 3439 1859 3455
rect 1793 3405 1809 3439
rect 1843 3405 1859 3439
rect 1793 3389 1859 3405
rect 1796 3358 1856 3389
rect 1796 2527 1856 2558
rect 1793 2511 1859 2527
rect 1793 2477 1809 2511
rect 1843 2477 1859 2511
rect 1793 2461 1859 2477
rect 2672 3514 2738 3530
rect 2672 3480 2688 3514
rect 2722 3480 2738 3514
rect 2672 3464 2738 3480
rect 2675 3433 2735 3464
rect 2675 2602 2735 2633
rect 2672 2586 2738 2602
rect 2672 2552 2688 2586
rect 2722 2552 2738 2586
rect 2672 2536 2738 2552
rect 3512 3501 3578 3517
rect 3512 3467 3528 3501
rect 3562 3467 3578 3501
rect 3512 3451 3578 3467
rect 3515 3420 3575 3451
rect 3515 2589 3575 2620
rect 3512 2573 3578 2589
rect 3512 2539 3528 2573
rect 3562 2539 3578 2573
rect 3512 2523 3578 2539
rect 946 1900 1036 1916
rect 946 1866 962 1900
rect 1020 1866 1036 1900
rect 946 1819 1036 1866
rect 946 972 1036 1019
rect 946 938 962 972
rect 1020 938 1036 972
rect 946 922 1036 938
rect 1806 1890 1896 1906
rect 1806 1856 1822 1890
rect 1880 1856 1896 1890
rect 1806 1809 1896 1856
rect 1806 962 1896 1009
rect 1806 928 1822 962
rect 1880 928 1896 962
rect 1806 912 1896 928
rect 2646 1910 2736 1926
rect 2646 1876 2662 1910
rect 2720 1876 2736 1910
rect 2646 1829 2736 1876
rect 2646 982 2736 1029
rect 2646 948 2662 982
rect 2720 948 2736 982
rect 2646 932 2736 948
rect 3466 1900 3556 1916
rect 3466 1866 3482 1900
rect 3540 1866 3556 1900
rect 3466 1819 3556 1866
rect 3466 972 3556 1019
rect 3466 938 3482 972
rect 3540 938 3556 972
rect 3466 922 3556 938
rect -4115 57 -4049 109
rect 953 639 1043 655
rect 953 605 969 639
rect 1027 605 1043 639
rect 953 567 1043 605
rect 953 129 1043 167
rect 953 95 969 129
rect 1027 95 1043 129
rect 953 79 1043 95
rect 1813 629 1903 645
rect 1813 595 1829 629
rect 1887 595 1903 629
rect 1813 557 1903 595
rect 1813 119 1903 157
rect 1813 85 1829 119
rect 1887 85 1903 119
rect 1813 69 1903 85
rect 2653 649 2743 665
rect 2653 615 2669 649
rect 2727 615 2743 649
rect 2653 577 2743 615
rect 2653 139 2743 177
rect 2653 105 2669 139
rect 2727 105 2743 139
rect 2653 89 2743 105
rect 3473 639 3563 655
rect 3473 605 3489 639
rect 3547 605 3563 639
rect 3473 567 3563 605
rect 3473 129 3563 167
rect 3473 95 3489 129
rect 3547 95 3563 129
rect 3473 79 3563 95
rect 973 -308 1039 -292
rect 973 -342 989 -308
rect 1023 -342 1039 -308
rect 973 -358 1039 -342
rect 976 -380 1036 -358
rect 976 -1202 1036 -1180
rect 973 -1218 1039 -1202
rect 973 -1252 989 -1218
rect 1023 -1252 1039 -1218
rect 973 -1268 1039 -1252
rect 1843 -288 1909 -272
rect 1843 -322 1859 -288
rect 1893 -322 1909 -288
rect 1843 -338 1909 -322
rect 1846 -360 1906 -338
rect 1846 -1182 1906 -1160
rect 1843 -1198 1909 -1182
rect 1843 -1232 1859 -1198
rect 1893 -1232 1909 -1198
rect 1843 -1248 1909 -1232
rect 2673 -298 2739 -282
rect 2673 -332 2689 -298
rect 2723 -332 2739 -298
rect 2673 -348 2739 -332
rect 2676 -370 2736 -348
rect 2676 -1192 2736 -1170
rect 2673 -1208 2739 -1192
rect 2673 -1242 2689 -1208
rect 2723 -1242 2739 -1208
rect 2673 -1258 2739 -1242
rect 3483 -278 3549 -262
rect 3483 -312 3499 -278
rect 3533 -312 3549 -278
rect 3483 -328 3549 -312
rect 3486 -350 3546 -328
rect 3486 -1172 3546 -1150
rect 3483 -1188 3549 -1172
rect 3483 -1222 3499 -1188
rect 3533 -1222 3549 -1188
rect 3483 -1238 3549 -1222
<< polycont >>
rect 969 3418 1003 3452
rect 969 2490 1003 2524
rect 1809 3405 1843 3439
rect 1809 2477 1843 2511
rect 2688 3480 2722 3514
rect 2688 2552 2722 2586
rect 3528 3467 3562 3501
rect 3528 2539 3562 2573
rect 962 1866 1020 1900
rect 962 938 1020 972
rect 1822 1856 1880 1890
rect 1822 928 1880 962
rect 2662 1876 2720 1910
rect 2662 948 2720 982
rect 3482 1866 3540 1900
rect 3482 938 3540 972
rect 969 605 1027 639
rect 969 95 1027 129
rect 1829 595 1887 629
rect 1829 85 1887 119
rect 2669 615 2727 649
rect 2669 105 2727 139
rect 3489 605 3547 639
rect 3489 95 3547 129
rect 989 -342 1023 -308
rect 989 -1252 1023 -1218
rect 1859 -322 1893 -288
rect 1859 -1232 1893 -1198
rect 2689 -332 2723 -298
rect 2689 -1242 2723 -1208
rect 3499 -312 3533 -278
rect 3499 -1222 3533 -1188
<< locali >>
rect 94 3957 221 3984
rect -992 3926 -865 3953
rect 918 3939 1072 3975
rect -2258 3577 -2108 3596
rect -2258 3502 -2251 3577
rect -2120 3502 -2108 3577
rect -2258 3293 -2108 3502
rect -992 3496 -865 3808
rect 94 3527 221 3839
rect 1059 3794 1072 3939
rect 1765 3930 1896 3957
rect 2594 3939 2752 3966
rect 3468 3939 3617 4002
rect 918 3554 1072 3794
rect 796 3520 892 3554
rect 1080 3520 1176 3554
rect 1765 3541 1896 3835
rect 2594 3616 2752 3844
rect 2515 3582 2611 3616
rect 2799 3582 2895 3616
rect 3468 3603 3617 3821
rect -856 3309 -716 3349
rect 230 3340 370 3380
rect -2158 3065 -2016 3116
rect 796 2422 830 3520
rect 953 3418 969 3452
rect 1003 3418 1019 3452
rect 1142 3375 1176 3520
rect 910 3359 944 3375
rect 1023 3359 1176 3375
rect 1023 3335 1028 3359
rect 910 2567 944 2583
rect 1062 3335 1176 3359
rect 1028 2567 1062 2583
rect 953 2490 969 2524
rect 1003 2490 1019 2524
rect 1142 2422 1176 3335
rect 796 2388 1176 2422
rect 1636 3507 1732 3541
rect 1920 3507 2016 3541
rect 1636 2409 1670 3507
rect 1765 3504 1896 3507
rect 1793 3405 1809 3439
rect 1843 3405 1859 3439
rect 1982 3362 2016 3507
rect 1750 3346 1784 3362
rect 1863 3346 2016 3362
rect 1863 3322 1868 3346
rect 1750 2554 1784 2570
rect 1902 3322 2016 3346
rect 1868 2554 1902 2570
rect 1793 2477 1809 2511
rect 1843 2477 1859 2511
rect 1982 2409 2016 3322
rect 2515 2484 2549 3582
rect 2594 3581 2752 3582
rect 2672 3480 2688 3514
rect 2722 3480 2738 3514
rect 2861 3437 2895 3582
rect 2629 3421 2663 3437
rect 2742 3421 2895 3437
rect 2742 3397 2747 3421
rect 2629 2629 2663 2645
rect 2781 3397 2895 3421
rect 2747 2629 2781 2645
rect 2672 2552 2688 2586
rect 2722 2552 2738 2586
rect 2861 2484 2895 3397
rect 2515 2450 2895 2484
rect 3355 3569 3451 3603
rect 3639 3569 3735 3603
rect 3355 2471 3389 3569
rect 3468 3559 3617 3569
rect 3512 3467 3528 3501
rect 3562 3467 3578 3501
rect 3701 3424 3735 3569
rect 3469 3408 3503 3424
rect 3582 3408 3735 3424
rect 3582 3384 3587 3408
rect 3469 2616 3503 2632
rect 3621 3384 3735 3408
rect 3587 2616 3621 2632
rect 3512 2539 3528 2573
rect 3562 2539 3578 2573
rect 3701 2471 3735 3384
rect 3355 2437 3735 2471
rect 4845 2666 4960 2690
rect 4845 2613 4857 2666
rect 4916 2613 4960 2666
rect 1636 2375 2016 2409
rect 4845 2168 4960 2613
rect 5805 2666 5922 2673
rect 5805 2618 5815 2666
rect 5896 2618 5922 2666
rect 5805 2133 5922 2618
rect 786 1968 1196 2002
rect 786 1906 820 1968
rect 946 1866 962 1900
rect 1020 1866 1036 1900
rect 900 1807 934 1823
rect 900 1015 934 1031
rect 1048 1807 1082 1823
rect 1048 1015 1082 1031
rect 946 938 962 972
rect 1020 938 1036 972
rect 786 870 820 932
rect 1162 870 1196 1968
rect 786 836 1196 870
rect 1646 1958 2056 1992
rect 1646 1896 1680 1958
rect 1806 1856 1822 1890
rect 1880 1856 1896 1890
rect 1760 1797 1794 1813
rect 1760 1005 1794 1021
rect 1908 1797 1942 1813
rect 1908 1005 1942 1021
rect 1806 928 1822 962
rect 1880 928 1896 962
rect 1646 860 1680 922
rect 2022 860 2056 1958
rect 1646 826 2056 860
rect 2486 1978 2896 2012
rect 2486 1916 2520 1978
rect 2646 1876 2662 1910
rect 2720 1876 2736 1910
rect 2600 1817 2634 1833
rect 2600 1025 2634 1041
rect 2748 1817 2782 1833
rect 2748 1025 2782 1041
rect 2646 948 2662 982
rect 2720 948 2736 982
rect 2486 880 2520 942
rect 2862 880 2896 1978
rect 2486 846 2896 880
rect 3306 1968 3716 2002
rect 3306 1906 3340 1968
rect 3466 1866 3482 1900
rect 3540 1866 3556 1900
rect 3420 1807 3454 1823
rect 3420 1015 3454 1031
rect 3568 1807 3602 1823
rect 3568 1015 3602 1031
rect 3466 938 3482 972
rect 3540 938 3556 972
rect 3306 870 3340 932
rect 3682 870 3716 1968
rect 3306 836 3716 870
rect 793 707 1203 741
rect 793 645 827 707
rect 953 605 969 639
rect 1027 605 1043 639
rect 907 555 941 571
rect 907 163 941 179
rect 1055 555 1089 571
rect 1055 163 1089 179
rect 953 95 969 129
rect 1027 95 1043 129
rect 793 27 827 89
rect 1169 27 1203 707
rect -2451 8 -2399 19
rect -2451 -26 -2446 8
rect -2412 -26 -2399 8
rect 793 -7 1203 27
rect 1653 697 2063 731
rect 1653 635 1687 697
rect 1813 595 1829 629
rect 1887 595 1903 629
rect 1767 545 1801 561
rect 1767 153 1801 169
rect 1915 545 1949 561
rect 1915 153 1949 169
rect 1813 85 1829 119
rect 1887 85 1903 119
rect 1653 17 1687 79
rect 2029 17 2063 697
rect 1653 -17 2063 17
rect 2493 717 2903 751
rect 2493 655 2527 717
rect 2653 615 2669 649
rect 2727 615 2743 649
rect 2607 565 2641 581
rect 2607 173 2641 189
rect 2755 565 2789 581
rect 2755 173 2789 189
rect 2653 105 2669 139
rect 2727 105 2743 139
rect 2493 37 2527 99
rect 2869 37 2903 717
rect 2493 3 2903 37
rect 3313 707 3723 741
rect 3313 645 3347 707
rect 3473 605 3489 639
rect 3547 605 3563 639
rect 3427 555 3461 571
rect 3427 163 3461 179
rect 3575 555 3609 571
rect 3575 163 3609 179
rect 3473 95 3489 129
rect 3547 95 3563 129
rect 3313 27 3347 89
rect 3689 27 3723 707
rect 4744 503 4845 506
rect 4738 471 4866 503
rect 5682 464 5795 521
rect 3313 -7 3723 27
rect -2451 -30 -2399 -26
rect 4846 -36 4907 249
rect 5801 -15 5882 247
rect 5873 -83 5882 -15
rect 5801 -85 5882 -83
rect 4846 -96 4907 -90
rect 816 -240 1196 -206
rect -2366 -1140 -2171 -1115
rect -2366 -1195 -2350 -1140
rect -2310 -1195 -2171 -1140
rect -879 -1126 -769 -1116
rect -879 -1156 -759 -1126
rect 260 -1130 370 -1120
rect 260 -1160 380 -1130
rect -2366 -1219 -2171 -1195
rect 816 -1320 850 -240
rect 973 -342 989 -308
rect 1023 -342 1039 -308
rect 930 -392 964 -376
rect 930 -1184 964 -1168
rect 1048 -392 1082 -376
rect 1162 -1090 1196 -240
rect 1082 -1140 1196 -1090
rect 1048 -1184 1082 -1168
rect 973 -1252 989 -1218
rect 1023 -1252 1039 -1218
rect 1162 -1320 1196 -1140
rect -1009 -1616 -889 -1336
rect -1009 -1666 -989 -1616
rect -999 -1686 -989 -1666
rect -919 -1666 -889 -1616
rect 130 -1620 250 -1340
rect 816 -1354 912 -1320
rect 1100 -1354 1196 -1320
rect 1686 -220 2066 -186
rect 1686 -1300 1720 -220
rect 1843 -322 1859 -288
rect 1893 -322 1909 -288
rect 1800 -372 1834 -356
rect 1800 -1164 1834 -1148
rect 1918 -372 1952 -356
rect 2032 -1060 2066 -220
rect 1952 -1100 2066 -1060
rect 1918 -1164 1952 -1148
rect 1843 -1232 1859 -1198
rect 1893 -1232 1909 -1198
rect 2032 -1300 2066 -1100
rect 1686 -1334 1782 -1300
rect 1970 -1334 2066 -1300
rect 2516 -230 2896 -196
rect 2516 -1310 2550 -230
rect 2673 -332 2689 -298
rect 2723 -332 2739 -298
rect 2630 -382 2664 -366
rect 2630 -1174 2664 -1158
rect 2748 -382 2782 -366
rect 2862 -1040 2896 -230
rect 2782 -1100 2896 -1040
rect 2748 -1174 2782 -1158
rect 2673 -1242 2689 -1208
rect 2723 -1242 2739 -1208
rect 2862 -1310 2896 -1100
rect -919 -1686 -909 -1666
rect 130 -1670 150 -1620
rect -999 -1696 -909 -1686
rect 140 -1690 150 -1670
rect 220 -1670 250 -1620
rect 980 -1630 1050 -1354
rect 220 -1690 230 -1670
rect 140 -1700 230 -1690
rect 1850 -1630 1940 -1334
rect 2516 -1344 2612 -1310
rect 2800 -1344 2896 -1310
rect 3326 -210 3706 -176
rect 3326 -1290 3360 -210
rect 3483 -312 3499 -278
rect 3533 -312 3549 -278
rect 3440 -362 3474 -346
rect 3440 -1154 3474 -1138
rect 3558 -362 3592 -346
rect 3672 -1040 3706 -210
rect 3592 -1110 3706 -1040
rect 3558 -1154 3592 -1138
rect 3483 -1222 3499 -1188
rect 3533 -1222 3549 -1188
rect 3672 -1290 3706 -1110
rect 3326 -1324 3422 -1290
rect 3610 -1324 3706 -1290
rect 1850 -1690 1870 -1630
rect 1930 -1690 1940 -1630
rect 2660 -1620 2780 -1344
rect 2660 -1680 2700 -1620
rect 1850 -1700 1940 -1690
rect 2750 -1680 2780 -1620
rect 3470 -1640 3570 -1324
rect 3470 -1710 3490 -1640
rect 3550 -1710 3570 -1640
rect 3470 -1720 3570 -1710
<< viali >>
rect -1001 3808 -820 3926
rect 85 3839 266 3957
rect -2251 3502 -2120 3577
rect 905 3794 1059 3939
rect 1711 3835 1919 3930
rect 2585 3844 2784 3939
rect 3454 3821 3653 3939
rect 969 3418 1003 3452
rect 910 2583 944 3359
rect 1028 2583 1062 3359
rect 969 2490 1003 2524
rect 1809 3405 1843 3439
rect 1750 2570 1784 3346
rect 1868 2570 1902 3346
rect 1809 2477 1843 2511
rect 2688 3480 2722 3514
rect 2629 2645 2663 3421
rect 2747 2645 2781 3421
rect 2688 2552 2722 2586
rect 3528 3467 3562 3501
rect 3469 2632 3503 3408
rect 3587 2632 3621 3408
rect 3528 2539 3562 2573
rect 4857 2613 4916 2666
rect 5815 2618 5896 2666
rect 962 1866 1020 1900
rect 900 1031 934 1807
rect 1048 1031 1082 1807
rect 962 938 1020 972
rect 1822 1856 1880 1890
rect 1760 1021 1794 1797
rect 1908 1021 1942 1797
rect 1822 928 1880 962
rect 2662 1876 2720 1910
rect 2600 1041 2634 1817
rect 2748 1041 2782 1817
rect 2662 948 2720 982
rect 3482 1866 3540 1900
rect 3420 1031 3454 1807
rect 3568 1031 3602 1807
rect 3482 938 3540 972
rect 969 605 1027 639
rect 907 179 941 555
rect 1055 179 1089 555
rect 969 95 1027 129
rect -2446 -26 -2412 8
rect 1829 595 1887 629
rect 1767 169 1801 545
rect 1915 169 1949 545
rect 1829 85 1887 119
rect 2669 615 2727 649
rect 2607 189 2641 565
rect 2755 189 2789 565
rect 2669 105 2727 139
rect 3489 605 3547 639
rect 3427 179 3461 555
rect 3575 179 3609 555
rect 3489 95 3547 129
rect 4837 -90 4912 -36
rect 5783 -83 5873 -15
rect -3854 -1213 -3816 -1176
rect -2350 -1195 -2310 -1140
rect 989 -342 1023 -308
rect 930 -1168 964 -392
rect 1048 -1168 1082 -392
rect 989 -1252 1023 -1218
rect -989 -1686 -919 -1616
rect 1859 -322 1893 -288
rect 1800 -1148 1834 -372
rect 1918 -1148 1952 -372
rect 1859 -1232 1893 -1198
rect 2689 -332 2723 -298
rect 2630 -1158 2664 -382
rect 2748 -1158 2782 -382
rect 2689 -1242 2723 -1208
rect 150 -1690 220 -1620
rect 970 -1700 1050 -1630
rect 3499 -312 3533 -278
rect 3440 -1138 3474 -362
rect 3558 -1138 3592 -362
rect 3499 -1222 3533 -1188
rect 1870 -1690 1930 -1630
rect 2700 -1700 2750 -1620
rect 3490 -1710 3550 -1640
<< metal1 >>
rect 3750 4029 5091 4035
rect -1856 3998 -1073 4000
rect -1856 3995 -617 3998
rect -1 3995 5091 4029
rect -1856 3957 5091 3995
rect -1856 3926 85 3957
rect -1856 3893 -1001 3926
rect -1867 3808 -1001 3893
rect -820 3839 85 3926
rect 266 3939 5091 3957
rect 266 3839 905 3939
rect -820 3808 905 3839
rect -1867 3794 905 3808
rect 1059 3930 2585 3939
rect 1059 3835 1711 3930
rect 1919 3844 2585 3930
rect 2784 3844 3454 3939
rect 1919 3835 3454 3844
rect 1059 3821 3454 3835
rect 3653 3821 5091 3939
rect 1059 3798 5091 3821
rect 1059 3794 5106 3798
rect -1867 3785 5106 3794
rect -1867 3763 52 3785
rect 3750 3773 5106 3785
rect -1867 3624 -1755 3763
rect -1087 3754 52 3763
rect -657 3751 52 3754
rect -2456 3577 -1755 3624
rect -2456 3502 -2251 3577
rect -2120 3502 -1755 3577
rect -2456 3480 -1755 3502
rect 2652 3514 2752 3527
rect 2652 3480 2688 3514
rect 2722 3480 2752 3514
rect -2456 3477 -1778 3480
rect -946 3379 -846 3439
rect 140 3410 240 3470
rect 2652 3467 2752 3480
rect 3492 3501 3592 3514
rect 3492 3467 3528 3501
rect 3562 3467 3592 3501
rect 933 3452 1033 3465
rect 3492 3454 3592 3467
rect 933 3418 969 3452
rect 1003 3418 1033 3452
rect 933 3405 1033 3418
rect 1773 3439 1873 3452
rect 1773 3405 1809 3439
rect 1843 3405 1873 3439
rect 1773 3392 1873 3405
rect 2623 3421 2669 3433
rect 904 3359 950 3371
rect -2237 3184 -2163 3230
rect -2309 2751 -2252 2762
rect -2309 2700 -2202 2751
rect -2309 2693 -2161 2700
rect -2309 2644 -2129 2693
rect -2272 2635 -2129 2644
rect -2242 2486 -2129 2635
rect 66 2653 143 2659
rect 904 2654 910 3359
rect -1020 2622 -943 2628
rect -1020 2568 -1012 2622
rect -954 2568 -943 2622
rect 66 2599 74 2653
rect 132 2599 143 2653
rect 66 2596 143 2599
rect 859 2648 910 2654
rect 74 2589 136 2596
rect 859 2594 867 2648
rect 859 2591 910 2594
rect 867 2584 910 2591
rect 904 2583 910 2584
rect 944 2583 950 3359
rect 904 2571 950 2583
rect 1022 3359 1068 3371
rect 1022 2583 1028 3359
rect 1062 2583 1068 3359
rect 1744 3346 1790 3358
rect 1744 2641 1750 3346
rect 1022 2571 1068 2583
rect 1699 2635 1750 2641
rect 1699 2581 1707 2635
rect 1699 2578 1750 2581
rect 1707 2571 1750 2578
rect -1020 2565 -943 2568
rect 1744 2570 1750 2571
rect 1784 2570 1790 3346
rect -1012 2558 -950 2565
rect 1744 2558 1790 2570
rect 1862 3346 1908 3358
rect 1862 2570 1868 3346
rect 1902 2570 1908 3346
rect 2623 2716 2629 3421
rect 2578 2710 2629 2716
rect 2578 2656 2586 2710
rect 2578 2653 2629 2656
rect 2586 2646 2629 2653
rect 2623 2645 2629 2646
rect 2663 2645 2669 3421
rect 2623 2633 2669 2645
rect 2741 3421 2787 3433
rect 2741 2645 2747 3421
rect 2781 2645 2787 3421
rect 3463 3408 3509 3420
rect 3463 2703 3469 3408
rect 2741 2633 2787 2645
rect 3418 2697 3469 2703
rect 3418 2643 3426 2697
rect 3418 2640 3469 2643
rect 3426 2633 3469 2640
rect 3463 2632 3469 2633
rect 3503 2632 3509 3408
rect 3463 2620 3509 2632
rect 3581 3408 3627 3420
rect 3581 2632 3587 3408
rect 3621 2632 3627 3408
rect 4821 2880 5106 3773
rect 4701 2843 5262 2880
rect 3581 2620 3627 2632
rect 4552 2666 6294 2843
rect 4552 2613 4857 2666
rect 4916 2618 5815 2666
rect 5896 2618 6294 2666
rect 4916 2613 6294 2618
rect 2672 2586 2742 2597
rect 2672 2583 2688 2586
rect 1862 2558 1908 2570
rect 2665 2552 2688 2583
rect 2722 2572 2742 2586
rect 3512 2573 3582 2584
rect 3512 2572 3528 2573
rect 2722 2552 3528 2572
rect 160 2516 230 2540
rect 2665 2539 3528 2552
rect 3562 2539 3582 2573
rect 953 2524 1023 2535
rect 953 2516 969 2524
rect -926 2496 -856 2509
rect 160 2496 969 2516
rect -926 2490 969 2496
rect 1003 2514 1023 2524
rect 2665 2534 3582 2539
rect 2665 2533 3574 2534
rect 2665 2523 3565 2533
rect 1793 2518 1863 2522
rect 2665 2518 2769 2523
rect 1793 2514 2769 2518
rect 1003 2511 2769 2514
rect 1003 2490 1809 2511
rect -926 2486 1809 2490
rect -2242 2477 1809 2486
rect 1843 2491 2769 2511
rect 4552 2501 6294 2613
rect 1843 2477 2727 2491
rect -2242 2432 2727 2477
rect -2242 2426 231 2432
rect -2227 2418 231 2426
rect 998 2424 2727 2432
rect 998 2423 1861 2424
rect -2227 2417 -878 2418
rect -1564 1985 -1498 2417
rect -4567 1983 -2450 1985
rect -2422 1983 -1498 1985
rect -4567 1882 -1498 1983
rect -4911 1825 -4809 1850
rect -4911 1773 -4883 1825
rect -4831 1773 -4809 1825
rect -4911 1755 -4809 1773
rect -4540 1705 -4491 1882
rect -4406 1825 -4336 1831
rect -4406 1824 -4396 1825
rect -4407 1823 -4396 1824
rect -4408 1773 -4396 1823
rect -4343 1773 -4336 1825
rect -4408 1767 -4336 1773
rect -4406 1765 -4336 1767
rect -4128 1822 -4026 1847
rect -4128 1770 -4100 1822
rect -4048 1770 -4026 1822
rect -4128 1752 -4026 1770
rect -3949 1713 -3900 1882
rect -3824 1820 -3722 1845
rect -3824 1768 -3796 1820
rect -3744 1768 -3722 1820
rect -3824 1750 -3722 1768
rect -3534 1815 -3432 1840
rect -3534 1763 -3506 1815
rect -3454 1763 -3432 1815
rect -3534 1745 -3432 1763
rect -3353 1705 -3313 1882
rect -3232 1813 -3130 1838
rect -3232 1761 -3204 1813
rect -3152 1761 -3130 1813
rect -3232 1743 -3130 1761
rect -2929 1815 -2827 1840
rect -2929 1763 -2901 1815
rect -2849 1763 -2827 1815
rect -2929 1745 -2827 1763
rect -2754 1703 -2718 1882
rect -2454 1880 -2393 1882
rect -2615 1822 -2513 1840
rect -2621 1815 -2513 1822
rect -2311 1820 -2209 1844
rect -2621 1770 -2587 1815
rect -2615 1763 -2587 1770
rect -2535 1763 -2513 1815
rect -2324 1819 -2209 1820
rect -2324 1772 -2283 1819
rect -2615 1745 -2513 1763
rect -2311 1767 -2283 1772
rect -2231 1767 -2209 1819
rect -2311 1749 -2209 1767
rect -2166 1704 -2120 1882
rect -2048 1817 -1946 1842
rect -2048 1765 -2020 1817
rect -1968 1765 -1946 1817
rect -2048 1747 -1946 1765
rect -1749 1811 -1647 1836
rect -1749 1759 -1721 1811
rect -1669 1759 -1647 1811
rect -1749 1741 -1647 1759
rect -1564 1745 -1498 1882
rect -1565 1703 -1498 1745
rect -130 2150 4000 2190
rect -130 780 -80 2150
rect 2650 1910 2732 1916
rect 950 1900 1032 1906
rect 950 1866 962 1900
rect 1020 1866 1032 1900
rect 950 1860 1032 1866
rect 1810 1890 1892 1896
rect 1810 1856 1822 1890
rect 1880 1856 1892 1890
rect 2650 1876 2662 1910
rect 2720 1876 2732 1910
rect 2650 1870 2732 1876
rect 3470 1900 3552 1906
rect 3470 1866 3482 1900
rect 3540 1866 3552 1900
rect 3470 1860 3552 1866
rect 1810 1850 1892 1856
rect 2558 1829 2633 1830
rect 2558 1824 2640 1829
rect 52 1814 118 1822
rect 52 1810 60 1814
rect 50 1760 60 1810
rect 113 1810 118 1814
rect 841 1819 931 1820
rect 841 1814 940 1819
rect 113 1760 120 1810
rect 50 1750 120 1760
rect 841 1760 864 1814
rect 923 1807 940 1814
rect 841 1750 900 1760
rect 240 1230 540 1270
rect 150 780 220 960
rect -130 740 220 780
rect 150 600 220 740
rect 480 790 540 1230
rect 894 1031 900 1750
rect 934 1031 940 1807
rect 894 1019 940 1031
rect 1042 1807 1088 1819
rect 1042 1031 1048 1807
rect 1082 1280 1088 1807
rect 1681 1809 1795 1819
rect 1681 1798 1800 1809
rect 1681 1739 1712 1798
rect 1765 1797 1800 1798
rect 1681 1727 1760 1739
rect 1082 1240 1350 1280
rect 1082 1031 1088 1240
rect 1042 1019 1088 1031
rect 950 972 1032 978
rect 950 938 962 972
rect 1020 938 1032 972
rect 950 932 1032 938
rect 960 790 1030 932
rect 480 750 1030 790
rect 480 430 540 750
rect 960 645 1030 750
rect 1290 780 1350 1240
rect 1754 1021 1760 1727
rect 1794 1021 1800 1797
rect 1754 1009 1800 1021
rect 1902 1797 1948 1809
rect 1902 1021 1908 1797
rect 1942 1270 1948 1797
rect 2558 1769 2568 1824
rect 2624 1817 2640 1824
rect 2558 1761 2600 1769
rect 1942 1230 2210 1270
rect 1942 1021 1948 1230
rect 1902 1009 1948 1021
rect 1810 962 1892 968
rect 1810 928 1822 962
rect 1880 928 1892 962
rect 1810 922 1892 928
rect 1820 780 1890 922
rect 1290 740 1890 780
rect 957 639 1039 645
rect 957 605 969 639
rect 1027 605 1039 639
rect 957 599 1039 605
rect 240 350 540 430
rect 901 555 947 567
rect 901 220 907 555
rect -4408 61 -4342 113
rect -4243 0 -4211 170
rect -4115 57 -4049 109
rect -3807 60 -3741 112
rect -3648 0 -3611 175
rect -3507 57 -3441 109
rect -3211 57 -3145 109
rect -3053 0 -3012 180
rect 40 170 130 210
rect 870 190 907 220
rect 850 179 907 190
rect 941 179 947 555
rect -2911 59 -2845 111
rect -2612 55 -2546 107
rect -2457 19 -2413 167
rect -2318 58 -2252 110
rect -2018 59 -1952 111
rect -2457 8 -2399 19
rect -2457 0 -2446 8
rect -4249 -26 -2446 0
rect -2412 0 -2399 8
rect -1862 0 -1814 154
rect -1723 56 -1657 108
rect -2412 -26 -1509 0
rect -4249 -34 -1509 -26
rect -4159 -1154 -4062 -34
rect -3648 -35 -3611 -34
rect -3053 -35 -3012 -34
rect -987 -295 -909 -276
rect -987 -297 -967 -295
rect -987 -319 -977 -297
rect -1028 -332 -977 -319
rect -1030 -339 -977 -332
rect -1039 -351 -977 -339
rect -911 -348 -909 -295
rect -912 -351 -909 -348
rect -1039 -357 -909 -351
rect -1039 -391 -965 -357
rect 40 -370 100 170
rect 850 167 947 179
rect 1049 555 1095 567
rect 1049 179 1055 555
rect 1089 440 1095 555
rect 1290 440 1350 740
rect 1820 635 1890 740
rect 2150 800 2210 1230
rect 2594 1041 2600 1761
rect 2634 1041 2640 1817
rect 2594 1029 2640 1041
rect 2742 1817 2788 1829
rect 2742 1041 2748 1817
rect 2782 1290 2788 1817
rect 3414 1812 3460 1819
rect 3367 1807 3460 1812
rect 3367 1803 3420 1807
rect 3367 1749 3392 1803
rect 3367 1740 3420 1749
rect 2782 1250 3050 1290
rect 2782 1041 2788 1250
rect 2742 1029 2788 1041
rect 2650 982 2732 988
rect 2650 948 2662 982
rect 2720 948 2732 982
rect 2650 942 2732 948
rect 2660 800 2730 942
rect 2150 760 2730 800
rect 1817 629 1899 635
rect 1817 595 1829 629
rect 1887 595 1899 629
rect 1817 589 1899 595
rect 1089 360 1350 440
rect 1761 545 1807 557
rect 1089 179 1095 360
rect 1761 200 1767 545
rect 1049 167 1095 179
rect 1720 169 1767 200
rect 1801 169 1807 545
rect 159 -289 241 -286
rect 159 -354 174 -289
rect 227 -354 241 -289
rect 159 -361 241 -354
rect 850 -360 910 167
rect 1720 157 1807 169
rect 1909 545 1955 557
rect 1909 169 1915 545
rect 1949 430 1955 545
rect 2150 430 2210 760
rect 2660 655 2730 760
rect 2990 790 3050 1250
rect 3414 1031 3420 1740
rect 3454 1031 3460 1807
rect 3414 1019 3460 1031
rect 3562 1807 3608 1819
rect 3562 1031 3568 1807
rect 3602 1280 3608 1807
rect 3602 1240 3870 1280
rect 3602 1031 3608 1240
rect 3562 1019 3608 1031
rect 3470 972 3552 978
rect 3470 938 3482 972
rect 3540 938 3552 972
rect 3470 932 3552 938
rect 3480 790 3550 932
rect 2990 750 3550 790
rect 2657 649 2739 655
rect 2657 615 2669 649
rect 2727 615 2739 649
rect 2657 609 2739 615
rect 1949 350 2210 430
rect 2601 565 2647 577
rect 1949 169 1955 350
rect 2601 230 2607 565
rect 1909 157 1955 169
rect 2550 189 2607 230
rect 2641 189 2647 565
rect 2550 177 2647 189
rect 2749 565 2795 577
rect 2749 189 2755 565
rect 2789 450 2795 565
rect 2990 450 3050 750
rect 3480 645 3550 750
rect 3810 920 3870 1240
rect 3940 920 4000 2150
rect 4853 2053 4931 2102
rect 5797 2023 5873 2073
rect 4926 1270 5195 1335
rect 4857 1118 4935 1172
rect 3810 919 4000 920
rect 4861 919 4921 1118
rect 3810 870 4921 919
rect 3477 639 3559 645
rect 3477 605 3489 639
rect 3547 605 3559 639
rect 3477 599 3559 605
rect 2789 370 3050 450
rect 3421 555 3467 567
rect 2789 189 2795 370
rect 3421 280 3427 555
rect 2749 177 2795 189
rect 3360 179 3427 280
rect 3461 179 3467 555
rect 957 129 1039 135
rect 957 95 969 129
rect 1027 95 1039 129
rect 957 89 1039 95
rect 971 -290 1052 -275
rect 971 -300 980 -290
rect 970 -343 980 -300
rect 1034 -343 1052 -290
rect 970 -350 1052 -343
rect 971 -351 1052 -350
rect 1720 -340 1780 157
rect 1817 119 1899 125
rect 1817 85 1829 119
rect 1887 85 1899 119
rect 1817 79 1899 85
rect 1841 -272 1934 -259
rect 1841 -280 1850 -272
rect 1840 -324 1850 -280
rect 1910 -324 1934 -272
rect 1840 -328 1934 -324
rect 1840 -330 1910 -328
rect 1720 -360 1810 -340
rect 2550 -350 2610 177
rect 3360 167 3467 179
rect 3569 555 3615 567
rect 3569 179 3575 555
rect 3609 440 3615 555
rect 3810 440 3870 870
rect 3922 867 4921 870
rect 4861 637 4921 867
rect 5126 928 5190 1270
rect 5873 1213 6126 1269
rect 5797 1095 5873 1145
rect 5805 928 5863 1095
rect 5126 855 5863 928
rect 6082 904 6124 1213
rect 5126 562 5190 855
rect 5805 686 5863 855
rect 6081 835 6276 904
rect 5795 633 5867 686
rect 4932 527 5190 562
rect 6082 523 6124 835
rect 5875 478 6124 523
rect 6082 477 6124 478
rect 3609 360 3870 440
rect 3609 179 3615 360
rect 4861 320 4930 375
rect 5801 320 5878 369
rect 3569 167 3615 179
rect 3360 150 3450 167
rect 2657 139 2739 145
rect 2657 105 2669 139
rect 2727 105 2739 139
rect 2657 99 2739 105
rect 2669 -283 2741 -270
rect 2669 -337 2682 -283
rect 2734 -337 2741 -283
rect 2669 -341 2741 -337
rect 3360 -330 3420 150
rect 3477 129 3559 135
rect 3477 95 3489 129
rect 3547 95 3559 129
rect 3477 89 3559 95
rect 4585 10 4765 14
rect 4585 -15 6002 10
rect 4585 -36 5783 -15
rect 4585 -90 4837 -36
rect 4912 -83 5783 -36
rect 5873 -83 6002 -15
rect 4912 -90 6002 -83
rect 4585 -105 6002 -90
rect 3477 -257 3549 -244
rect 3477 -310 3486 -257
rect 3539 -270 3549 -257
rect 3539 -310 3550 -270
rect 3477 -312 3499 -310
rect 3533 -312 3550 -310
rect 3477 -317 3550 -312
rect 3480 -320 3550 -317
rect 3360 -350 3450 -330
rect -1039 -455 -982 -391
rect 40 -460 130 -370
rect 850 -380 940 -360
rect 1720 -372 1840 -360
rect 850 -392 970 -380
rect 850 -450 930 -392
rect -2363 -1118 -1865 -1116
rect -2369 -1140 -1823 -1118
rect -4159 -1176 -3796 -1154
rect -4159 -1213 -3854 -1176
rect -3816 -1213 -3796 -1176
rect -4159 -1239 -3796 -1213
rect -2369 -1195 -2350 -1140
rect -2310 -1195 -1823 -1140
rect 924 -1168 930 -450
rect 964 -1168 970 -392
rect 924 -1180 970 -1168
rect 1042 -392 1088 -380
rect 1042 -1168 1048 -392
rect 1082 -1168 1088 -392
rect 1720 -430 1800 -372
rect 1794 -1148 1800 -430
rect 1834 -1148 1840 -372
rect 1794 -1160 1840 -1148
rect 1912 -372 1958 -360
rect 1912 -1148 1918 -372
rect 1952 -1148 1958 -372
rect 2550 -370 2640 -350
rect 3360 -362 3480 -350
rect 2550 -382 2670 -370
rect 2550 -440 2630 -382
rect 1912 -1160 1958 -1148
rect 2624 -1158 2630 -440
rect 2664 -1158 2670 -382
rect 1042 -1180 1088 -1168
rect 2624 -1170 2670 -1158
rect 2742 -382 2788 -370
rect 2742 -1158 2748 -382
rect 2782 -1158 2788 -382
rect 3360 -420 3440 -362
rect 3434 -1138 3440 -420
rect 3474 -1138 3480 -362
rect 3434 -1150 3480 -1138
rect 3552 -362 3598 -350
rect 3552 -1138 3558 -362
rect 3592 -1138 3598 -362
rect 3552 -1150 3598 -1138
rect 3908 -627 4160 -616
rect 4585 -627 4765 -105
rect 3908 -742 4765 -627
rect 2742 -1170 2788 -1158
rect 3470 -1188 3560 -1180
rect -2369 -1219 -1823 -1195
rect 1830 -1198 1920 -1190
rect -2369 -1222 -2294 -1219
rect -4159 -1247 -4062 -1239
rect -1969 -1594 -1823 -1219
rect -989 -1266 -899 -1216
rect 960 -1218 1050 -1210
rect 150 -1270 240 -1220
rect 960 -1252 989 -1218
rect 1023 -1252 1050 -1218
rect 1830 -1232 1859 -1198
rect 1893 -1232 1920 -1198
rect 1830 -1240 1920 -1232
rect 2660 -1208 2750 -1200
rect 2660 -1242 2689 -1208
rect 2723 -1242 2750 -1208
rect 3470 -1222 3499 -1188
rect 3533 -1222 3560 -1188
rect 3470 -1230 3560 -1222
rect 2660 -1250 2750 -1242
rect 960 -1260 1050 -1252
rect -1969 -1596 -1206 -1594
rect -1969 -1598 -645 -1596
rect -1969 -1600 -65 -1598
rect 3908 -1600 4160 -742
rect 4585 -753 4765 -742
rect -1969 -1616 4160 -1600
rect -1969 -1686 -989 -1616
rect -919 -1620 4160 -1616
rect -919 -1686 150 -1620
rect -1969 -1690 150 -1686
rect 220 -1630 2700 -1620
rect 220 -1690 970 -1630
rect -1969 -1700 970 -1690
rect 1050 -1690 1870 -1630
rect 1930 -1690 2700 -1630
rect 1050 -1700 2700 -1690
rect 2750 -1640 4160 -1620
rect 2750 -1700 3490 -1640
rect -1969 -1710 3490 -1700
rect 3550 -1656 4160 -1640
rect 3550 -1710 4062 -1656
rect -1969 -1722 4062 -1710
rect -1941 -1726 4062 -1722
rect -1941 -1730 -1206 -1726
rect -677 -1730 4062 -1726
rect -677 -1731 -65 -1730
rect 3768 -1747 4062 -1730
<< via1 >>
rect -1012 2568 -954 2622
rect 74 2599 132 2653
rect 867 2594 910 2648
rect 910 2594 925 2648
rect 1707 2581 1750 2635
rect 1750 2581 1765 2635
rect 2586 2656 2629 2710
rect 2629 2656 2644 2710
rect 3426 2643 3469 2697
rect 3469 2643 3484 2697
rect -4883 1773 -4831 1825
rect -4396 1773 -4343 1825
rect -4100 1770 -4048 1822
rect -3796 1768 -3744 1820
rect -3506 1763 -3454 1815
rect -3204 1761 -3152 1813
rect -2901 1763 -2849 1815
rect -2587 1763 -2535 1815
rect -2283 1767 -2231 1819
rect -2020 1765 -1968 1817
rect -1721 1759 -1669 1811
rect 60 1760 113 1814
rect 864 1807 923 1814
rect 864 1760 900 1807
rect 900 1760 923 1807
rect 1712 1797 1765 1798
rect 1712 1739 1760 1797
rect 1760 1739 1765 1797
rect 2568 1817 2624 1824
rect 2568 1769 2600 1817
rect 2600 1769 2624 1817
rect -967 -297 -911 -295
rect -977 -348 -911 -297
rect -977 -351 -912 -348
rect 3392 1749 3420 1803
rect 3420 1749 3448 1803
rect 174 -354 227 -289
rect 980 -308 1034 -290
rect 980 -342 989 -308
rect 989 -342 1023 -308
rect 1023 -342 1034 -308
rect 980 -343 1034 -342
rect 1850 -288 1910 -272
rect 1850 -322 1859 -288
rect 1859 -322 1893 -288
rect 1893 -322 1910 -288
rect 1850 -324 1910 -322
rect 2682 -298 2734 -283
rect 2682 -332 2689 -298
rect 2689 -332 2723 -298
rect 2723 -332 2734 -298
rect 2682 -337 2734 -332
rect 3486 -278 3539 -257
rect 3486 -310 3499 -278
rect 3499 -310 3533 -278
rect 3533 -310 3539 -278
<< metal2 >>
rect 2578 2710 2655 2716
rect 2578 2677 2586 2710
rect 66 2653 143 2659
rect 2562 2656 2586 2677
rect 2644 2656 2655 2710
rect 3418 2697 3495 2703
rect 3418 2664 3426 2697
rect -1020 2622 -943 2628
rect -1020 2589 -1012 2622
rect -1036 2568 -1012 2589
rect -954 2568 -943 2622
rect 66 2620 74 2653
rect -1036 2565 -943 2568
rect 50 2599 74 2620
rect 132 2599 143 2653
rect 859 2648 936 2654
rect 859 2615 867 2648
rect 50 2596 143 2599
rect 50 2590 140 2596
rect 843 2594 867 2615
rect 925 2594 936 2648
rect 2562 2653 2655 2656
rect 2562 2647 2652 2653
rect 2562 2646 2648 2647
rect 1699 2635 1776 2641
rect 1699 2602 1707 2635
rect 843 2591 936 2594
rect 50 2589 136 2590
rect -1036 2559 -946 2565
rect -1036 2558 -950 2559
rect -1036 2275 -996 2558
rect -1037 2253 -996 2275
rect -4911 1842 -4809 1850
rect -4128 1842 -4026 1847
rect -3824 1842 -3722 1845
rect -2311 1842 -2209 1844
rect -4911 1836 -1660 1842
rect -4911 1825 -1647 1836
rect -4911 1773 -4883 1825
rect -4831 1787 -4396 1825
rect -4831 1773 -4809 1787
rect -4911 1755 -4809 1773
rect -4408 1773 -4396 1787
rect -4343 1822 -1647 1825
rect -4343 1787 -4100 1822
rect -4343 1773 -4336 1787
rect -4408 1767 -4336 1773
rect -4406 1765 -4336 1767
rect -4128 1770 -4100 1787
rect -4048 1820 -1647 1822
rect -4048 1787 -3796 1820
rect -4048 1770 -4026 1787
rect -4128 1752 -4026 1770
rect -3824 1768 -3796 1787
rect -3744 1819 -1647 1820
rect -3744 1815 -2283 1819
rect -3744 1787 -3506 1815
rect -3744 1768 -3722 1787
rect -3824 1750 -3722 1768
rect -3534 1763 -3506 1787
rect -3454 1813 -2901 1815
rect -3454 1787 -3204 1813
rect -3454 1763 -3432 1787
rect -3534 1745 -3432 1763
rect -3232 1761 -3204 1787
rect -3152 1787 -2901 1813
rect -3152 1761 -3130 1787
rect -3232 1743 -3130 1761
rect -2929 1763 -2901 1787
rect -2849 1787 -2587 1815
rect -2849 1763 -2827 1787
rect -2929 1745 -2827 1763
rect -2615 1763 -2587 1787
rect -2535 1787 -2283 1815
rect -2535 1763 -2513 1787
rect -2615 1745 -2513 1763
rect -2311 1767 -2283 1787
rect -2231 1817 -1647 1819
rect -2231 1787 -2020 1817
rect -2231 1767 -2209 1787
rect -2311 1749 -2209 1767
rect -2048 1765 -2020 1787
rect -1968 1811 -1647 1817
rect -1968 1787 -1721 1811
rect -1968 1765 -1946 1787
rect -2048 1747 -1946 1765
rect -1749 1759 -1721 1787
rect -1669 1759 -1647 1811
rect -1749 1741 -1647 1759
rect -1037 -184 -997 2253
rect 50 1821 90 2589
rect 843 2585 933 2591
rect 843 2584 929 2585
rect 843 2318 883 2584
rect 840 2309 883 2318
rect 1683 2581 1707 2602
rect 1765 2581 1776 2635
rect 1683 2578 1776 2581
rect 1683 2572 1773 2578
rect 1683 2571 1769 2572
rect 1683 2311 1723 2571
rect 2562 2379 2602 2646
rect 3402 2643 3426 2664
rect 3484 2643 3495 2697
rect 3402 2640 3495 2643
rect 3402 2634 3492 2640
rect 3402 2633 3488 2634
rect 3402 2381 3442 2633
rect 2558 2371 2602 2379
rect 50 1814 120 1821
rect 50 1760 60 1814
rect 113 1760 120 1814
rect 840 1820 879 2309
rect 840 1814 931 1820
rect 1682 1819 1725 2311
rect 2558 1830 2599 2371
rect 3399 2358 3442 2381
rect 2558 1824 2633 1830
rect 840 1776 864 1814
rect 50 1750 120 1760
rect 841 1760 864 1776
rect 923 1760 931 1814
rect 841 1750 931 1760
rect 1681 1798 1795 1819
rect 1681 1739 1712 1798
rect 1765 1739 1795 1798
rect 2558 1769 2568 1824
rect 2624 1769 2633 1824
rect 3399 1813 3440 2358
rect 3380 1812 3442 1813
rect 2558 1761 2633 1769
rect 3367 1803 3448 1812
rect 3367 1749 3392 1803
rect 3367 1740 3448 1749
rect 1681 1727 1795 1739
rect -1037 -248 -906 -184
rect -992 -276 -910 -248
rect 3267 -257 3551 -231
rect 1841 -260 1934 -259
rect 3267 -260 3486 -257
rect 1050 -268 1719 -267
rect 1841 -268 3486 -260
rect 1050 -272 3486 -268
rect -992 -280 -909 -276
rect -992 -281 -147 -280
rect -992 -282 240 -281
rect 1050 -282 1850 -272
rect -992 -289 1850 -282
rect -992 -295 174 -289
rect -992 -297 -967 -295
rect -992 -304 -977 -297
rect -987 -351 -977 -304
rect -911 -341 174 -295
rect -911 -348 -909 -341
rect -171 -344 174 -341
rect -912 -351 -909 -348
rect -987 -357 -909 -351
rect 159 -354 174 -344
rect 227 -290 1850 -289
rect 227 -343 980 -290
rect 1034 -324 1850 -290
rect 1910 -283 3486 -272
rect 1910 -324 2682 -283
rect 1034 -337 2682 -324
rect 2734 -310 3486 -283
rect 3539 -310 3551 -257
rect 2734 -318 3551 -310
rect 2734 -337 3311 -318
rect 1034 -338 3311 -337
rect 1034 -343 1719 -338
rect 1908 -341 3311 -338
rect 227 -354 1719 -343
rect 2659 -342 3311 -341
rect 2659 -349 2741 -342
rect 159 -357 1719 -354
rect 159 -358 1054 -357
rect 159 -361 241 -358
use sky130_fd_pr__nfet_01v8_BLLLZK  sky130_fd_pr__nfet_01v8_BLLLZK_0
timestamp 1702646674
transform 1 0 -943 0 1 -786
box -226 -610 226 610
use sky130_fd_pr__nfet_01v8_BLLLZK  sky130_fd_pr__nfet_01v8_BLLLZK_1
timestamp 1702646674
transform 1 0 196 0 1 -790
box -226 -610 226 610
use sky130_fd_pr__nfet_01v8_MMDDFP  sky130_fd_pr__nfet_01v8_MMDDFP_0
timestamp 1702652280
transform 1 0 -3033 0 1 940
box -1657 -1010 1657 1010
use sky130_fd_pr__nfet_01v8_MVKWCS  sky130_fd_pr__nfet_01v8_MVKWCS_0
timestamp 1702646674
transform 1 0 188 0 1 357
box -241 -410 241 410
use sky130_fd_pr__nfet_01v8_RB2QBJ  sky130_fd_pr__nfet_01v8_RB2QBJ_0
timestamp 1702648458
transform 1 0 5835 0 1 505
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_RB2QBJ  sky130_fd_pr__nfet_01v8_RB2QBJ_1
timestamp 1702648458
transform 1 0 4896 0 1 505
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_9K6AJ9  sky130_fd_pr__pfet_01v8_9K6AJ9_0
timestamp 1702648458
transform 1 0 5836 0 1 1584
box -211 -619 211 619
use sky130_fd_pr__pfet_01v8_9K6AJ9  sky130_fd_pr__pfet_01v8_9K6AJ9_1
timestamp 1702648458
transform 1 0 4893 0 1 1608
box -211 -619 211 619
use sky130_fd_pr__pfet_01v8_882MTD  sky130_fd_pr__pfet_01v8_882MTD_0
timestamp 1702652280
transform 1 0 -2201 0 1 2941
box -226 -419 226 419
use sky130_fd_pr__pfet_01v8_AYYC2A  sky130_fd_pr__pfet_01v8_AYYC2A_0
timestamp 1702646674
transform 1 0 181 0 1 1409
box -241 -619 241 619
use sky130_fd_pr__pfet_01v8_YSNZTD  sky130_fd_pr__pfet_01v8_YSNZTD_0
timestamp 1702647685
transform 1 0 -893 0 1 2945
box -226 -619 226 619
use sky130_fd_pr__pfet_01v8_YSNZTD  sky130_fd_pr__pfet_01v8_YSNZTD_1
timestamp 1702647685
transform 1 0 193 0 1 2976
box -226 -619 226 619
use sky130_fd_pr__res_xhigh_po_0p35_9HMPAT  sky130_fd_pr__res_xhigh_po_0p35_9HMPAT_0
timestamp 1702652280
transform 1 0 -3083 0 1 -1113
box -948 -484 948 484
<< labels >>
rlabel via1 -4877 1777 -4836 1821 1 Vctrl
port 1 n
rlabel metal1 -2432 3528 -2358 3579 1 Vdd
port 2 n
rlabel metal1 -1683 -1696 -1609 -1645 1 GND
port 3 n
rlabel metal1 6175 846 6249 897 1 Vout
port 4 n
<< end >>
